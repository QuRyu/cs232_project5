library ieee;
library ieee.std_logic_1164.all;

entity ROM is 
    port (
        addr : std_logic_vector (3 downto 0);
        data : std_logic_vector (9 downto 0)
    );
end entity;

architecture rlt of ROM is 

begin

end rlt;
